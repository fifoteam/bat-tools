//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : chk_flhide
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/27 13:52:31	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module chk_flhide # (
	parameter	DATA_WIDTH		= 8		,	//����λ��
	parameter	CHANNEL_NUM		= 4		,	//ͨ����
	parameter	STOP_ON_ERROR	= 1			//���ִ���ʱ�Ƿ�ֹͣ
	)
	(
	input										clk			,	//ʱ��
	input										i_fval		,	//����Ч
	input										i_lval		,	//����Ч
	input	[DATA_WIDTH*CHANNEL_NUM-1:0]		iv_pix_data		//����Ч
	);

	//	ref signals


	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	����fval=0ʱ���������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!i_fval) begin
			if(i_lval==1'b1 || iv_pix_data!={(DATA_WIDTH*CHANNEL_NUM){1'b0}}) begin
				$display("%m: at time %t ERROR: when fval=0,lval pix_data not 0", $time);
				if(STOP_ON_ERROR==1) begin
					$stop;
				end
			end
		end
	end

	//	-------------------------------------------------------------------------------------
	//	����fval=0ʱ���������
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!i_lval) begin
			if(iv_pix_data!={(DATA_WIDTH*CHANNEL_NUM){1'b0}}) begin
				$display("%m: at time %t ERROR: when lval=0,pix_data not 0", $time);
				if(STOP_ON_ERROR==1) begin
					$stop;
				end
			end
		end
	end

endmodule
