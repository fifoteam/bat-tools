//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : chipscope_top
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/10/27 10:21:13	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module chipscope_top (
	input				CLK			,
	input	[16:0]		TRIG0		,
	output	[15:0]		ASYNC_OUT
	);

	//	ref signals
	wire	[35:0]			CONTROL0	;
	wire	[35:0]			CONTROL1	;

	//	ref ARCHITECTURE
	chipscope_icon_user1_2port chipscope_icon_user1_2port_inst (
	.CONTROL0	(CONTROL0	),
	.CONTROL1	(CONTROL1	)
	);

	chipscope_ila_w17_d1k chipscope_ila_w17_d1k_inst (
	.CONTROL	(CONTROL0	),
	.CLK		(CLK		),
	.TRIG0		(TRIG0		)
	);

	chipscope_vio_16_async_out chipscope_vio_16_async_out_inst (
	.CONTROL	(CONTROL1	),
	.ASYNC_OUT	(ASYNC_OUT	)
	);


endmodule
