//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : chk_data_align
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/3/19 13:48:24	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
//`timescale 1ns/1ps
`timescale 1ns/1ns
//-------------------------------------------------------------------------------------------------

module chk_data_align # (
	parameter		REG_WD					= 32	,	//�Ĵ���λ��
	parameter		DATA_DEPTH 				= 64	,	//�������
	parameter		DATA_IN_WIDTH			= 10	,	//��������λ��
	parameter		DATA_OUT_WIDTH			= 32	,	//�������λ��
	parameter		STOP_ON_ERROR			= 1			//���ִ����Ƿ�ֹͣ
	)
	(
	input							i_chk_en		,	//��鿪��
	input	[REG_WD-1:0]			iv_pixel_format	,	//���ظ�ʽ�Ĵ�����0x01080001:Mono8��0x01100003:Mono10��0x01080008:BayerGR8��0x0110000C:BayerGR10
	input							clk_in			,	//����ʱ��
	input							i_fval_in		,	//���볡�ź�
	input							i_lval_in		,	//�������ź�
	input	[DATA_IN_WIDTH-1:0]		iv_pix_data_in	,	//��������
	input							clk_out			,	//���ʱ��
	input							i_fval_out		,	//������ź�
	input							i_lval_out		,	//������ź�
	input	[DATA_OUT_WIDTH-1:0]	iv_pix_data_out		//�������

	);

	//	ref signals
	reg		[DATA_IN_WIDTH-1:0]		mem	[DATA_DEPTH-1:0]	;
	reg		[11:0]					addr_a	= 12'b0	;	//��ַ12bit����������4k
	reg		[11:0]					addr_b	= 12'b0	;
	reg								format8_sel	= 1'b0	;
	wire	[DATA_OUT_WIDTH-1:0]	data_group_8	;
	wire	[DATA_OUT_WIDTH-1:0]	data_group_10	;

	//	ref ARCHITECTURE

	//  ===============================================================================================
	//	ref ***�ж����ݸ�ʽ***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	Mono8		- 0x01080001	-> 0x1081	-> 0001,0000,1000,,,,0001
	//	Mono10		- 0x01100003	-> 0x1103	-> 0001,0001,0000,,,,0011
	//	BayerGR8	- 0x01080008	-> 0x1088	-> 0001,0000,1000,,,,1000
	//	BayerGR10	- 0x0110000C	-> 0x110C	-> 0001,0001,0000,,,,1100
	//											   --------!-!-------!!!!
	//                                                     ^    ^       ^------bit0
	//                                             bit20---|    |---bit16
	//	����� ! �ģ����ǲ���Ƚϵ�bit.�ֱ��� bit
	//  -------------------------------------------------------------------------------------
	//  -------------------------------------------------------------------------------------
	//	format8_sel
	//	1.�ж����ظ�ʽ�Ƿ�ѡ��8bit���ظ�ʽ
	//	2.ʹ��6bit�ж�����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk_out) begin
		case({iv_pixel_format[20],iv_pixel_format[19],iv_pixel_format[3:0]})
			6'b010001	: format8_sel	<= 1'b1;
			6'b011000	: format8_sel	<= 1'b1;
			default		: format8_sel	<= 1'b0;
		endcase
	end

	//  ===============================================================================================
	//	ref ***�洢������***
	//  ===============================================================================================
	//  -------------------------------------------------------------------------------------
	//	����ʱ����
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk_in) begin
		if(i_fval_in==1'b1 && i_lval_in==1'b1 && i_chk_en==1'b1) begin
			addr_a	<= addr_a + 1'b1;
		end
	end

	always @ (posedge clk_in) begin
		if(i_fval_in==1'b1 && i_lval_in==1'b1 && i_chk_en==1'b1) begin
			mem[addr_a]	<= iv_pix_data_in;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	���ʱ����
	//	1.���ظ�ʽ��8bit��ÿ�����ڣ���ַ+4
	//	1.���ظ�ʽ��10bit��ÿ�����ڣ���ַ+2
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk_out) begin
		if(i_fval_out==1'b1 && i_lval_out==1'b1 && i_chk_en==1'b1) begin
			if(format8_sel) begin
				addr_b	<= addr_b + 3'b100;
			end
			else begin
				addr_b	<= addr_b + 2'b10;
			end
		end
	end

	//	-------------------------------------------------------------------------------------
	//	�������
	//	1.��������ź�ʹ���ұȽϿ��ش�ʱ�����ܱȽϣ�����û���κζ���
	//	2.��������������ram�е����ݲ�һ�������ӡ������Ϣ�����ݲ�����ѡ���Ƿ�ֹͣ��
	//	-------------------------------------------------------------------------------------
	assign	data_group_8	= {mem[addr_b+3][DATA_IN_WIDTH-1:DATA_IN_WIDTH-8],mem[addr_b+2][DATA_IN_WIDTH-1:DATA_IN_WIDTH-8],mem[addr_b+1][DATA_IN_WIDTH-1:DATA_IN_WIDTH-8],mem[addr_b][DATA_IN_WIDTH-1:DATA_IN_WIDTH-8]};
	assign	data_group_10	= {6'b0,mem[addr_b+1],6'b0,mem[addr_b]};
	always @ (posedge clk_out) begin
		if(i_fval_out==1'b1 && i_lval_out==1'b1 && i_chk_en==1'b1) begin
			if(format8_sel) begin
				if(iv_pix_data_out!=data_group_8) begin
					$display ("%m:time is %t ERROR input data is %h,mem data is %h",$time,iv_pix_data_out,data_group_8);
					if(STOP_ON_ERROR) begin
						$stop;
					end
				end
			end
			else begin
				if(iv_pix_data_out!=data_group_10) begin
					$display ("%m:time is %t ERROR input data is %h,mem data is %h",$time,iv_pix_data_out,data_group_10);
					if(STOP_ON_ERROR) begin
						$stop;
					end
				end
			end

		end
	end






endmodule
