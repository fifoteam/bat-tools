//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : bfm_encrypt
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/10 15:46:57	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------
`define		TESTCASE	testcase1
module bfm_encrypt ();

	//	ref signals
	reg			i_encrypt_state		= 1'b0;

	//	ref ARCHITECTURE

	//	-------------------------------------------------------------------------------------
	//	--ref ����
	//	-------------------------------------------------------------------------------------
	//	-------------------------------------------------------------------------------------
	//	����״̬
	//	-------------------------------------------------------------------------------------
	task encrypt_low;
		begin
			#1
			i_encrypt_state	= 1'b0;
		end
	endtask

	task encrypt_high;
		begin
			#1
			i_encrypt_state	= 1'b1;
		end
	endtask



endmodule
