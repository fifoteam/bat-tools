//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : chk_pulse_width
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2015/4/14 10:41:05	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :
//              1)  : ... ...
//
//              2)  : ... ...
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module chk_pulse_width # (
	parameter		LARGE1_SMALL0		= 0		,	//1-���ڵ��ڸ������ȣ�0-С�ڵ��ڸ�������
	parameter		PULSE_POL			= 1		,	//���弫�ԣ�1-�ߵ�ƽ��0-�͵�ƽ
	parameter		COUNT_WIDHT			= 16	,	//���������Ŀ��
	parameter		STOP_ON_ERROR		= 1			//���ִ����Ƿ�ֹͣ
	)
	(
	input						clk				,	//ʱ��
	input						i_chk_en		,	//��⿪��
	input						i_din			,	//�����ź�
	input	[COUNT_WIDHT-1:0]	iv_pulse_width	,	//������
	output						o_error			//�����źţ���ʾ���ִ���ֱ��ʹ�ܹرղŻ�����
	);

	//	ref signals

	//FSM Parameter Define
	parameter	S_IDLE		= 1'd0;
	parameter	S_PULSE		= 1'd1;

	reg		[0:0]	current_state	= S_IDLE;
	reg		[0:0]	next_state		= S_IDLE;

	//FSM for sim
	// synthesis translate_off
	reg		[63:0]			state_ascii;
	always @ ( * ) begin
		case(current_state)
			1'd0 :	state_ascii	<= "S_IDLE";
			1'd1 :	state_ascii	<= "S_PULSE";
		endcase
	end
	// synthesis translate_on

	reg		[2:0]				din_shift	= 3'b000;
	wire						din_rise	;
	wire						din_fall	;
	wire						first_edge	;
	wire						second_edge	;
	reg		[COUNT_WIDHT-1:0]	pulse_width_cnt	= {COUNT_WIDHT{1'b0}};
	reg							error_reg	= 1'b0;

	//	ref ARCHITECTURE

	//	===============================================================================================
	//	ref ***��ʱ ȡ����***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	�������ź�ȡ����
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		din_shift	<= {din_shift[1:0],i_din};
	end
	assign	din_rise	= (din_shift[2:1]==2'b01) ? 1'b1 : 1'b0;
	assign	din_fall	= (din_shift[2:1]==2'b10) ? 1'b1 : 1'b0;

	//	-------------------------------------------------------------------------------------
	//	����ǵ����壬���һ���������½��أ��ڶ���������������
	//	����Ǹ����壬���һ�������������أ��ڶ����������½���
	//	-------------------------------------------------------------------------------------
	assign	first_edge	= (PULSE_POL==0 && din_fall==1'b1) ? 1'b1 : ((PULSE_POL==1 && din_rise==1'b1) ? 1'b1 : 1'b0);
	assign	second_edge	= (PULSE_POL==0 && din_rise==1'b1) ? 1'b1 : ((PULSE_POL==1 && din_fall==1'b1) ? 1'b1 : 1'b0);

	//	===============================================================================================
	//	ref ***�ж�����***
	//	===============================================================================================
	//	-------------------------------------------------------------------------------------
	//	���������
	//	-------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(current_state==S_IDLE) begin
			pulse_width_cnt	<= {COUNT_WIDHT{1'b0}};
		end
		else begin
			pulse_width_cnt	<= pulse_width_cnt + 1'b1;
		end
	end

	//	-------------------------------------------------------------------------------------
	//	�����ź�
	//	1.ֻ�е�����ź�ȡ����ʱ�򣬲�������
	//	2.�����ڼ���״̬���ҵڶ����½��ص���ʱ���ж�����
	//	-------------------------------------------------------------------------------------
	generate
		//	-------------------------------------------------------------------------------------
		//	��������
		//	-------------------------------------------------------------------------------------
		if(LARGE1_SMALL0==1) begin
			always @ (posedge clk) begin
				if(!i_chk_en) begin
					error_reg	<= 1'b0;
				end
				if(current_state==S_PULSE && second_edge==1'b1) begin
					if(pulse_width_cnt+1 >= iv_pulse_width) begin
						error_reg	<= 1'b1;
					end
				end
			end
		end
		//	-------------------------------------------------------------------------------------
		//	���խ����
		//	-------------------------------------------------------------------------------------
		else begin
			always @ (posedge clk) begin
				if(!i_chk_en) begin
					error_reg	<= 1'b0;
				end
				if(current_state==S_PULSE && second_edge==1'b1) begin
					if(pulse_width_cnt+1 <= iv_pulse_width) begin
						error_reg	<= 1'b1;
					end
				end
			end
		end
	endgenerate
	assign	o_error	= error_reg;

	//	-------------------------------------------------------------------------------------
	//	������
	//	-------------------------------------------------------------------------------------
	always @ (posedge error_reg) begin
		$display("%m: at time %t ERROR: pulse width check", $time);
		if(STOP_ON_ERROR) begin
			$stop;
		end
	end

	//	===============================================================================================
	//	ref ***״̬��***
	//	===============================================================================================
	//FSM Sequential Logic
	always @ (posedge clk) begin
		if(!i_chk_en) begin
			current_state	<= S_IDLE;
		end else begin
			current_state	<= next_state;
		end
	end

	//FSM Conbinatial Logic
	always @ ( * ) begin
		case(current_state)
			//	-------------------------------------------------------------------------------------
			//	�������źŵĵ�һ�����ص���ʱ����ʼ����
			//	-------------------------------------------------------------------------------------
			S_IDLE	:
			if(first_edge) begin
				next_state	= S_PULSE;
			end
			else begin
				next_state	= S_IDLE;
			end
			//	-------------------------------------------------------------------------------------
			//	�������źŵĵڶ������ص���ʱ��ֹͣ����
			//	-------------------------------------------------------------------------------------
			S_PULSE	:
			if(second_edge) begin
				next_state	= S_IDLE;
			end
			else begin
				next_state	= S_PULSE;
			end
			default	:
			next_state	= S_IDLE;
		endcase
	end





endmodule
